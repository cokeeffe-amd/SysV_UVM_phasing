// Forward declarations to resolve circular dependencies
//not sure what this does but CoPilot insists on it
typedef class my_phase_base;
typedef class PhaseScheduler;
