`ifndef PHASE_TYPES_SV
    `define PHASE_TYPES_SV

    // Forward declarations to resolve circular dependencies
    // NB: code does not work without these!
    typedef class my_phase_base;
    typedef class PhaseScheduler;

`endif // PHASE_TYPES_SV
